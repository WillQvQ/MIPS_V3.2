`timescale 1ns / 1ps

module mem#(parameter N = 64, L = 128)(
    input   logic           clk, 
    input   logic           dword,
    input   logic           memread,
    input   logic [1:0]     memwrite,
    input   logic [N-1:0]   dataadr, writedata,
    input   logic [31:0]    instradr,
    output  logic [31:0]    instr,
    output  logic [N-1:0]   readdata,
    input   logic [7:0]     checka,
    output  logic [31:0]    check,
    output  logic           ready,
    input   logic [7:0]     rx_data,
    output  logic [31:0]    rx_check,
    output  logic [31:0]    rx_checkh,
    output  logic [31:0]    rx_checkl
);
    logic [N-1:0] RAM [L-1:0];
    logic [31:0]  word;
    logic [N-1:0] rdata;
    logic [7:0]   cnt;
    initial ready = 1;
    initial cnt = 8'b0;
    initial $readmemh("C:/Users/will131/Documents/workspace/MIPS_V3.2/memfile.dat",RAM);
    assign instr = instradr[2] ? RAM[instradr[31:3]][31:0] : RAM[instradr[31:3]][63:32];
    assign rdata = dword ? RAM[dataadr[N-1:3]] : {32'b0,word};
    assign check = checka[0] ? RAM[checka[7:1]][31:0] : RAM[checka[7:1]][63:32];
    assign word = dataadr[2] ? RAM[dataadr[N-1:3]][31:0] : RAM[dataadr[N-1:3]][63:32];
    assign rx_check = rx_data[0] ? RAM[rx_data[7:1]][31:0] : RAM[rx_data[7:1]][63:32];
    assign rx_checkh = RAM[rx_data[7:1]][63:32];
    assign rx_checkl = RAM[rx_data[7:1]][31:0];
    always @(negedge clk)begin
        if((cnt==0) & memread)begin
            ready <= 0;
            cnt <= 8'd20;
        end
        else if (memwrite==2)begin
            case (dataadr[2:0])
                3'b111:  RAM[dataadr[N-1:3]][7:0]   <= writedata[7:0];
                3'b110:  RAM[dataadr[N-1:3]][15:8]  <= writedata[7:0];
                3'b101:  RAM[dataadr[N-1:3]][23:16] <= writedata[7:0];
                3'b100:  RAM[dataadr[N-1:3]][31:24] <= writedata[7:0];
                3'b011:  RAM[dataadr[N-1:3]][39:32] <= writedata[7:0];
                3'b010:  RAM[dataadr[N-1:3]][47:40] <= writedata[7:0];
                3'b001:  RAM[dataadr[N-1:3]][55:48] <= writedata[7:0];
                3'b000:  RAM[dataadr[N-1:3]][63:56] <= writedata[7:0];
            endcase
            ready <= 0;
            cnt <= 8'd20;
        end
        else if (memwrite==1)begin
            case (dataadr[2])
                0:  RAM[dataadr[N-1:3]][63:32]  <= writedata[31:0];
                1:  RAM[dataadr[N-1:3]][31:0]   <= writedata[31:0];
            endcase
            ready <= 0;
            cnt <= 8'd20;
        end
        if (memwrite==3)begin
            RAM[dataadr[N-1:3]] <= writedata;
            ready <= 0;
            cnt <= 8'd20;
        end
        else if(cnt!=0)begin
            if(cnt==1)begin
                readdata <= rdata;
                ready <= 1;
                cnt <= 0;
            end
            else cnt <= cnt - 1;
        end
    end 
endmodule